
module alt_clk_div (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
